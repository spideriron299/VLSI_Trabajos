LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY mux IS
	PORT(SEL : IN INTEGER RANGE 0 TO 3;
	        CP: OUT INTEGER RANGE 0 TO 9);
			  
END ENTITY;

ARCHITECTURE BEAS OF mux IS
BEGIN

	
	WITH SEL SELECT
		  CP <= 9 WHEN 0,
				  5 WHEN 1, 
				  2 WHEN 2, 
				  0 WHEN OTHERS;

END BEAS;
